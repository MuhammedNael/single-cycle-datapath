module control(
    input conditionBalv,
    input conditionBgtzal,
    input [5:0] opcode,
    input [5:0] funcCode,
    output reg [1:0] RegDst,
    output reg ALUSrc,
    output reg MemToReg,
    output reg RegWrite,
    output reg MemRead,
    output reg MemWrite,
    output reg Branch,
    output reg [1:0] ALUOp,
    output reg [1:0] Jump,
    output reg Brnv,
    output reg Nandi,
    output reg MuxReg,
    output reg Balv,
    output reg Bgtzal,
    output reg Jrsal,
    output reg StatusRegWrite
);

    always @(*) begin
        // Default values
        RegDst = 2'b00;
        ALUSrc = 0;
        MemToReg = 0;
        RegWrite = 0;
        MemRead = 0;
        MemWrite = 0;
        Branch = 0;
        ALUOp = 2'b00;
        Jump = 2'b00;
        Brnv = 0;
        Nandi = 0;
        MuxReg = 0;
        Balv = 0;
        Bgtzal = 0;
        Jrsal = 0;
        StatusRegWrite = 0;

        case (opcode)
            6'b000000: begin // R-format
                case (funcCode)
                    6'b100111: begin // Jmnor (R - F)
                        RegDst = 2'b10;
                        ALUSrc = 0;
                        MemToReg = 0;
                        RegWrite = 1;
                        MemRead = 0;
                        MemWrite = 0;
                        Branch = 0;
                        ALUOp = 2'b10;
                        Jump = 2'b11;
                        Brnv = 0;
                        Nandi = 0;
                        MuxReg = 0;
                        Balv = 0;
                        Bgtzal = 0;
                        Jrsal = 0;
                        StatusRegWrite = 0;
                    end
                    6'b010101: begin // Brnv (R - F)
                        RegDst = 2'b00;
                        ALUSrc = 0;
                        MemToReg = 0;
                        RegWrite = 0;
                        MemRead = 0;
                        MemWrite = 0;
                        Branch = 0;
                        ALUOp = 2'b10;
                        Jump = 2'b01;
                        Brnv = 1;
                        Nandi = 0;
                        MuxReg = 0;
                        Balv = 0;
                        Bgtzal = 0;
                        Jrsal = 0;
                        StatusRegWrite = 0;
                    end
                    default: begin
                        RegDst = 2'b01;
                        ALUSrc = 0;
                        MemToReg = 0;
                        RegWrite = 1;
                        MemRead = 0;
                        MemWrite = 0;
                        Branch = 0;
                        ALUOp = 2'b10;
                        Jump = 2'b01;
                        Brnv = 0;
                        Nandi = 0;
                        MuxReg = 1;
                        Balv = 0;
                        Bgtzal = 0;
                        Jrsal = 0;
                        StatusRegWrite = 1;
                    end
                endcase
            end

            6'b100011: begin // lw
                RegDst = 2'b00;
                ALUSrc = 1;
                MemToReg = 1;
                RegWrite = 1;
                MemRead = 1;
                MemWrite = 0;
                Branch = 0;
                ALUOp = 2'b00;
                Jump = 2'b01;
                Brnv = 0;
                Nandi = 0;
                MuxReg = 1;
                Balv = 0;
                Bgtzal = 0;
                Jrsal = 0;
                StatusRegWrite = 0;
            end
            6'b101011: begin // sw
                RegDst = 2'b00;
                ALUSrc = 1;
                MemToReg = 0;
                RegWrite = 0;
                MemRead = 0;
                MemWrite = 1;
                Branch = 0;
                ALUOp = 2'b00;
                Jump = 2'b01;
                Brnv = 0;
                Nandi = 0;
                MuxReg = 0;
                Balv = 0;
                Bgtzal = 0;
                Jrsal = 0;
                StatusRegWrite = 0;
            end
            6'b000100: begin // beq
                RegDst = 2'b00;
                ALUSrc = 0;
                MemToReg = 0;
                RegWrite = 0;
                MemRead = 0;
                MemWrite = 0;
                Branch = 1;
                ALUOp = 2'b01;
                Jump = 2'b01;
                Brnv = 0;
                Nandi = 0;
                MuxReg = 0;
                Balv = 0;
                Bgtzal = 0;
                Jrsal = 0;
                StatusRegWrite = 0;
            end
            6'b010000: begin // Nandi
                RegDst = 2'b00;
                ALUSrc = 1;
                MemToReg = 0;
                RegWrite = 1;
                MemRead = 0;
                MemWrite = 0;
                Branch = 0;
                ALUOp = 2'b11;
                Jump = 2'b01;
                Brnv = 0;
                Nandi = 1;
                MuxReg = 1;
                Balv = 0;
                Bgtzal = 0;
                Jrsal = 0;
                StatusRegWrite = 1;
            end
            6'b100001: begin // Bgtzal
                RegDst = 2'b11;
                ALUSrc = 0;
                MemToReg = 0;
                RegWrite = conditionBgtzal;
                MemRead = 0;
                MemWrite = 0;
                Branch = 0;
                ALUOp = 2'b00;
                Jump = 2'b00;
                Brnv = 0;
                Nandi = 0;
                MuxReg = 0;
                Balv = 0;
                Bgtzal = 1;
                Jrsal = 0;
                StatusRegWrite = 0;
            end
            6'b100000: begin // Balv
                RegDst = 2'b10;
                ALUSrc = 0;
                MemToReg = 0;
                RegWrite = conditionBalv;
                MemRead = 0;
                MemWrite = 0;
                Branch = 0;
                ALUOp = 2'b00;
                Jump = 2'b00;
                Brnv = 0;
                Nandi = 0;
                MuxReg = 0;
                Balv = 1;
                Bgtzal = 0;
                Jrsal = 0;
                StatusRegWrite = 0;
            end
            6'b010001: begin // Jrsal
                RegDst = 2'b00;
                ALUSrc = 0;
                MemToReg = 1;
                RegWrite = 0;
                MemRead = 1;
                MemWrite = 1;
                Branch = 0;
                ALUOp = 2'b00;
                Jump = 2'b10;
                Brnv = 0;
                Nandi = 0;
                MuxReg = 0;
                Balv = 0;
                Bgtzal = 0;
                Jrsal = 1;
                StatusRegWrite = 0;
            end
        endcase
    end
endmodule

